// unsaved_tb.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module unsaved_tb (
	);

	wire        unsaved_inst_clk_bfm_clk_clk;                     // unsaved_inst_clk_bfm:clk -> [unsaved_inst:clk_clk, unsaved_inst_reset_bfm:clk]
	wire        unsaved_inst_video_vga_controller_conduits_blank; // unsaved_inst:video_vga_controller_conduits_BLANK -> unsaved_inst_video_vga_controller_conduits_bfm:sig_BLANK
	wire  [7:0] unsaved_inst_video_vga_controller_conduits_b;     // unsaved_inst:video_vga_controller_conduits_B -> unsaved_inst_video_vga_controller_conduits_bfm:sig_B
	wire  [7:0] unsaved_inst_video_vga_controller_conduits_r;     // unsaved_inst:video_vga_controller_conduits_R -> unsaved_inst_video_vga_controller_conduits_bfm:sig_R
	wire        unsaved_inst_video_vga_controller_conduits_clk;   // unsaved_inst:video_vga_controller_conduits_CLK -> unsaved_inst_video_vga_controller_conduits_bfm:sig_CLK
	wire  [7:0] unsaved_inst_video_vga_controller_conduits_g;     // unsaved_inst:video_vga_controller_conduits_G -> unsaved_inst_video_vga_controller_conduits_bfm:sig_G
	wire        unsaved_inst_video_vga_controller_conduits_hs;    // unsaved_inst:video_vga_controller_conduits_HS -> unsaved_inst_video_vga_controller_conduits_bfm:sig_HS
	wire        unsaved_inst_video_vga_controller_conduits_sync;  // unsaved_inst:video_vga_controller_conduits_SYNC -> unsaved_inst_video_vga_controller_conduits_bfm:sig_SYNC
	wire        unsaved_inst_video_vga_controller_conduits_vs;    // unsaved_inst:video_vga_controller_conduits_VS -> unsaved_inst_video_vga_controller_conduits_bfm:sig_VS
	wire        unsaved_inst_reset_bfm_reset_reset;               // unsaved_inst_reset_bfm:reset -> unsaved_inst:reset_reset_n

	unsaved unsaved_inst (
		.clk_clk                             (unsaved_inst_clk_bfm_clk_clk),                     //                           clk.clk
		.reset_reset_n                       (unsaved_inst_reset_bfm_reset_reset),               //                         reset.reset_n
		.video_vga_controller_conduits_CLK   (unsaved_inst_video_vga_controller_conduits_clk),   // video_vga_controller_conduits.CLK
		.video_vga_controller_conduits_HS    (unsaved_inst_video_vga_controller_conduits_hs),    //                              .HS
		.video_vga_controller_conduits_VS    (unsaved_inst_video_vga_controller_conduits_vs),    //                              .VS
		.video_vga_controller_conduits_BLANK (unsaved_inst_video_vga_controller_conduits_blank), //                              .BLANK
		.video_vga_controller_conduits_SYNC  (unsaved_inst_video_vga_controller_conduits_sync),  //                              .SYNC
		.video_vga_controller_conduits_R     (unsaved_inst_video_vga_controller_conduits_r),     //                              .R
		.video_vga_controller_conduits_G     (unsaved_inst_video_vga_controller_conduits_g),     //                              .G
		.video_vga_controller_conduits_B     (unsaved_inst_video_vga_controller_conduits_b)      //                              .B
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) unsaved_inst_clk_bfm (
		.clk (unsaved_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) unsaved_inst_reset_bfm (
		.reset (unsaved_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (unsaved_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm unsaved_inst_video_vga_controller_conduits_bfm (
		.sig_B     (unsaved_inst_video_vga_controller_conduits_b),     // conduit.B
		.sig_BLANK (unsaved_inst_video_vga_controller_conduits_blank), //        .BLANK
		.sig_CLK   (unsaved_inst_video_vga_controller_conduits_clk),   //        .CLK
		.sig_G     (unsaved_inst_video_vga_controller_conduits_g),     //        .G
		.sig_HS    (unsaved_inst_video_vga_controller_conduits_hs),    //        .HS
		.sig_R     (unsaved_inst_video_vga_controller_conduits_r),     //        .R
		.sig_SYNC  (unsaved_inst_video_vga_controller_conduits_sync),  //        .SYNC
		.sig_VS    (unsaved_inst_video_vga_controller_conduits_vs)     //        .VS
	);

endmodule
